library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity deneme is
port (
      -- inputs
      a : in std_logic;
      b : in std_logic; 
      -- outputs
      z : out std_logic
      );
end deneme;

architecture Behavioral of deneme is
    -- helper vars (wires and stuff as signal)
    
begin
    -- algorithm

end Behavioral;
